`timescale 1ns/1ps

module alu_test;


reg[31:0] i_datain,gr1,gr2;


wire[31:0] c;
wire[3:0] ALUCr;
wire[0:0] zero, overflow, neg;



alu testalu(i_datain, gr1, gr2, c, zero, overflow, neg);

initial
begin

$display("--------------------------------------------------------------------");
$display("instruction:op:func:ALUCr:  gr1   :  gr2   :   c    : reg_a  : reg_b");
$display("--------------------------------------------------------------------");
$monitor("   %h:%h: %h :  %h  :%h:%h:%h:%h:%h",
testalu.i_dataIn, testalu.op, testalu.func, testalu.ALUCr, gr1, gr2, c, testalu.reg_a, testalu.reg_b);


/*//// 		R type instructions test 		////*/

//// logical left shift

#10 $display("   <<< sll >>>");
	i_datain<= 32'b0000_0000_0000_0001_0001_0000_0100_0000;
	gr2<= 32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<= 32'b0000_0000_0000_0001_0001_0000_1000_0000;
	gr2<= 32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<= 32'b0000_0000_0000_0001_0001_0000_0100_0000;
	gr2<= 32'b0100_0000_0100_0000_0100_0000_0100_0000;

#10 i_datain<= 32'b0000_0000_0000_0001_0001_0001_0000_0000;
	gr2<= 32'b0100_0000_0100_0000_0100_0000_0100_0000;


//// sllv

#10 $display("   <<< sllv >>>");
	i_datain <= 32'b0000_0000_0000_0001_0001_000000_000100;
	gr1 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0001_0000;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_000000_000100;
	gr1 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_000000_000100;
	gr1 <= 32'b0100_0000_0100_0000_0100_0000_0100_0000;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_000000_000100;
	gr1 <= 32'b0100_0000_0100_0000_0100_0000_0100_0000;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;

//// logical right shift

#10 $display("   <<< srl >>>");
	i_datain <= 32'b000000_00000_00001_00010_00010_000010;
	gr2 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain <= 32'b000000_00000_00001_00010_01000_000010;
	gr2 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain <= 32'b000000_00000_00001_00010_00010_000010;
	gr2 <= 32'b1111_1111_1111_1111_1111_1111_1101_1101;

#10 i_datain <= 32'b000000_00000_00001_00010_01000_000010;
	gr2 <= 32'b1111_1111_1111_1111_1111_1111_1101_1101;

//// srlv

#10 $display("   <<< srlv >>>");
	i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0110;
	gr1 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0110;
	gr1 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0110;
	gr1 <= 32'b0101_0101_0101_0101_0101_0101_0101_0101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0110;
	gr1 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;


//// sra

#10 $display("   <<< sra >>>");
	i_datain <= 32'b0000_0000_0000_0001_0001_0000_1000_0011;
	gr2 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0010_0000_0011;
	gr2 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0000_1000_0011;
	gr2 <= 32'b0101_0101_0101_0101_0101_0101_0101_0101;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0010_0000_0011;
	gr2 <= 32'b0101_0101_0101_0101_0101_0101_0101_0101;


//// srav
	
#10 $display("   <<< srav >>>");
	i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0111;
	gr1 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0111;
	gr1 <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0111;
	gr1 <= 32'b0101_0101_0101_0101_0101_0101_0101_0101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;

#10 i_datain <= 32'b0000_0000_0000_0001_0001_0000_0000_0111;
	gr1 <= 32'b0101_0101_0101_0101_0101_0101_0101_0101;
	gr2 <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;


//// add

#10 $display("   <<< add >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100000;
	gr1 <= 32'b000000_11010_01010_11101_10101_100000;
	gr2 <= 32'b101001_10101_10101_10010_11111_101001;

#10 i_datain <= 32'b000000_00000_00001_00010_00000_100000;
	gr1 <= 32'b100000_11010_01010_11101_10101_100000;
	gr2 <= 32'b101001_10101_10101_10010_11111_101001;


//// addu

#10	$display("   <<< addu >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100001;
	gr1 <= 32'b000000_11010_01010_11101_10101_100000;
	gr2 <= 32'b101001_10101_10101_10010_11111_101001;

#10 i_datain <= 32'b000000_00000_00001_00010_00000_100001;
	gr1 <= 32'b100000_11010_01010_11101_10101_100000;
	gr2 <= 32'b101001_10101_10101_10010_11111_101001;

//// sub

#10	$display("   <<< sub >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100010;
	gr1 <= 32'b000101_10101_01010_00101_00000_111011;
	gr2 <= 32'b100100_10010_11010_10010_00000_101101;

#10 i_datain <= 32'b000000_00000_00001_00010_00000_100010;
	gr1 <= 32'b010101_10101_01010_00101_00000_111011;
	gr2 <= 32'b110100_10010_11010_10010_00000_101101;

//// subu
	
#10	$display("   <<< subu >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100011;
	gr1 <= 32'b000101_10101_01010_00101_00000_111011;
	gr2 <= 32'b100100_10010_11010_10010_00000_101101;

#10	i_datain <= 32'b000000_00000_00001_00010_00000_100011;
	gr1 <= 32'b010101_10101_01010_00101_00000_111011;
	gr2 <= 32'b110100_10010_11010_10010_00000_101101;

//// mult

#10	$display("   <<< mult >>>");
	i_datain <= 32'b000000_00100_01000_00000_00000_011000;
	gr1 <= 32'b000100_10000_10100_10101_01100_101010;
	gr2 <= 32'b111010_10100_10100_10100_10101_101010;

#10 i_datain <= 32'b000000_00100_01000_00000_00000_011000;
	gr1 <= 32'b100100_10000_10100_10101_01100_101010;
	gr2 <= 32'b111010_10100_10100_10100_10101_101010;

//// multu

#10	$display("   <<< multu >>>");
	i_datain <= 32'b000000_00100_01000_00000_00000_011001;
	gr1 <= 32'b000100_10000_10100_10101_01100_101010;
	gr2 <= 32'b111010_10100_10100_10100_10101_101010;


#10 i_datain <= 32'b000000_00100_01000_00000_00000_011001;
	gr1 <= 32'b100100_10000_10100_10101_01100_101010;
	gr2 <= 32'b111010_10100_10100_10100_10101_101010;

//// div

#10	$display("   <<< div >>>");
	i_datain <= 32'b000000_00100_01000_00000_00000_011010;
	gr1 <= 32'b010010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

#10 i_datain <= 32'b000000_00100_01000_00000_00000_011010;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

//// divu
	
#10	$display("   <<< divu >>>");
	i_datain <= 32'b000000_00100_01000_00000_00000_011011;
	gr1 <= 32'b010010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

#10 i_datain <= 32'b000000_00100_01000_00000_00000_011011;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

//// and

#10	$display("   <<< and >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100100;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

#10 i_datain <= 32'b000000_00000_00001_00010_00000_100100;
	gr1 <= 32'b000010_10100_10010_10101_10101_111001;
	gr2 <= 32'b000101_11111_11000_10011_10000_101001;

//// nor

#10	$display("   <<< nor >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100111;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

#10 i_datain <= 32'b000000_00000_00001_00010_00000_100111;
	gr1 <= 32'b000010_10100_10010_10101_10101_111001;
	gr2 <= 32'b000101_11111_11000_10011_10000_101001;

//// or

#10	$display("   <<< or >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100101;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

#10 i_datain <= 32'b000000_00000_00001_00010_00000_100101;
	gr1 <= 32'b000010_10100_10010_10101_10101_111001;
	gr2 <= 32'b000101_11111_11000_10011_10000_101001;


//// xor

#10	$display("   <<< xor >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_100110;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

#10 i_datain <= 32'b000000_00000_00001_00010_00000_100110;
	gr1 <= 32'b000010_10100_10010_10101_10101_111001;
	gr2 <= 32'b000101_11111_11000_10011_10000_101001;


//// slt

#10	$display("   <<< slt >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_101010;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;

//// sltu

#10	$display("   <<< sltu >>>");
	i_datain <= 32'b000000_00000_00001_00010_00000_101011;
	gr1 <= 32'b111010_10100_10010_10101_10101_111111;
	gr2 <= 32'b000001_10101_11101_10011_11010_101001;


/*//// 		I type instructions test 		////*/

//// addi

#10 $display("   <<< addi >>>");
	i_datain <= 32'b001000_00000_10001_10010_00000_100000;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;

//// addiu

#10 $display("   <<< addiu >>>");
	i_datain <= 32'b001001_00000_10001_10010_00000_100000;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;

//// andi

#10 $display("   <<< andi >>>");
	i_datain <= 32'b001100_00000_00001_01010_10010_101010;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;

//// ori

#10 $display("   <<< ori >>>");
	i_datain <= 32'b001101_00000_00001_01010_00000_110101;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;

//// xori

#10 $display("   <<< xori >>>");
	i_datain <= 32'b001110_00000_00001_01010_00000_110101;
	gr1 <= 32'b110010_10100_10010_10101_10101_111111;

//// slti

#10 $display("   <<< slti >>>");
	i_datain <= 32'b001010_00000_00001_00100_00010_001010;
	gr1 <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;

//// sltiu

#10 $display("   <<< sltiu >>>");
	i_datain <= 32'b001011_00000_00001_10100_00010_001010;
	gr1 <= 32'b0000_0000_0000_0000_0100_0000_0000_1111;

//// beq

#10 $display("   <<< beq >>>");
	i_datain <= 32'b000100_00000_00001_00001_10000_011111;
	gr1 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;
	gr2 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;

#10 i_datain <= 32'b000100_00000_00001_00001_10000_011111;
	gr1 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;
	gr2 <= 32'b0000_0000_1010_1111_1010_1101_1000_1000;

//// bne

#10 $display("   <<< bne >>>");
	i_datain <= 32'b000101_00000_00001_00001_10000_011111;
	gr1 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;
	gr2 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;

#10 i_datain <= 32'b000101_00000_00001_00001_10000_011111;
	gr1 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;
	gr2 <= 32'b0000_0000_1010_1111_1010_1101_1000_1000;

//// lw

#10 $display("   <<< lw >>>");
	i_datain <= 32'b100011_00000_00001_00010_10101_101010;
	gr1 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;

//// sw

#10 $display("   <<< sw >>>");
	i_datain <= 32'b101011_00000_00001_00010_10101_101010;
	gr1 <= 32'b0000_0000_1010_1111_1010_1101_1000_0000;



#10 $finish;
end

endmodule